`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   23:41:14 06/22/2018
// Design Name:   count
// Module Name:   C:/Users/magnifico/Desktop/FPGA/Huffman/Huffman/count_test.v
// Project Name:  Huffman
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: count
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module count_test;

	// Inputs
	reg CLK;
	reg nRST;
	reg input_over;
	reg [1023:0] CHARACTER_IN;

	// Outputs
	wire [129:0] FREQUENT_OUT;
	wire count_over;

	// Instantiate the Unit Under Test (UUT)
	count uut (
		.CLK(CLK), 
		.nRST(nRST), 
		.input_over(input_over),
		.CHARACTER_IN(CHARACTER_IN), 
		.FREQUENT_OUT(FREQUENT_OUT),
		.count_over(count_over)
	);

	initial begin
		// Initialize Inputs
		CLK = 0;
		nRST = 0;
		input_over = 1'b1;
		CHARACTER_IN = 1024'b1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_0010_0011_0011_0100_0100_0100_0101_0101_0101_0101_0110_0110_0110_0110_0110_0111_0111_0111_0111_0111_0111_1000_1000_1000_1000_1000_1000_1000_1001_1001_1001_1001_1001_1001_1001_1001;

		// Wait 100 ns for global reset to finish
		#100;
     nRST = 1;
		// Add stimulus here

	end
	parameter DELAY = 1;
	always 
		#DELAY CLK = ~ CLK;
      
endmodule

