`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:59:59 06/21/2018
// Design Name:   main
// Module Name:   C:/Users/magnifico/Desktop/FPGA/Huffman/Huffman/main_test.v
// Project Name:  Huffman
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: main
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module main_test;

	// Inputs
	reg CLK;
	reg nRST;
	reg [3:0] input_data;
	reg input_start;

	// Outputs
	wire data;
	wire done;
	wire output_start;

	// Instantiate the Unit Under Test (UUT)
	main uut (
		.CLK(CLK), 
		.nRST(nRST),
		.input_data(input_data),
		.input_start(input_start),
		.data(data),
		.done(done),
		.output_start(output_start)
	);
	
	reg [1023:0] character;
	integer K;

	initial begin
		// Initialize Inputs
		CLK = 0;
		nRST = 0;
		character <= 1024'b1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_1001_1000_0111_0110_0101_0100_0011_0010_0001_0000_0010_0011_0011_0100_0100_0100_0101_0101_0101_0101_0110_0110_0110_0110_0110_0111_0111_0111_0111_0111_0111_1000_1000_1000_1000_1000_1000_1000_1001_1001_1001_1001_1001_1001_1001_1001;

		// Wait 100 ns for global reset to finish
		#100;
        
	nRST = 1;
	#5;
	input_start = 1;
	for (K = 0; K < 256; K = K + 1)
	begin
	  input_data[3:0] = character[3:0];
	  character = #2 {4'b0000,character[1023:4]};
	end
		// Add stimulus here

	end
	parameter DELAY = 1;
	always 
		#DELAY CLK = ~ CLK;

endmodule

